`ifndef APB_MASTER_STATES_VH
`define APB_MASTER_STATES_VH

// Define the states of the APB master
`define IDLE   2'b00  // Idle state
`define SETUP  2'b01  // Setup state
`define ACCESS 2'b10  // Access state

`endif // APB_MASTER_STATES_VH
